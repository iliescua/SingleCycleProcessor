library ieee;
use ieee.std_logic_1164.all;

entity bmux32bit is
port(D0,D1 : in std_logic_vector(31 downto 0);
	  S : in std_logic;
	  Y : out std_logic_vector(31 downto 0));
end entity bmux32bit;

architecture Dataflow of bmux32bit is 
begin

	with S select
		Y <= D0 when '0',
			  D1 when '1';
			  
end architecture Dataflow;