--Bmux2to1
--Andrew Iliescu
--4/29/18
library ieee;
use ieee.std_logic_1164.all;

entity bmux2to1 is--begin entity
port(D0,D1: in std_logic_vector(31 downto 0);
	  S : in std_logic;
	  Y : out std_logic_vector(31 downto 0));
end bmux2to1;--end entity

architecture Dataflow of bmux2to1 is--begin dataflow architecture
begin 

	with S select--with select picks the appropriate location based on selector bits
		Y <= D1 when '1',
			  D0 when '0';

end architecture Dataflow;--end dataflow architecture