--LR
--Andrew Iliescu
--4/29/18
library ieee;
use ieee.std_logic_1164.all;

entity lr is
port(input : in std_logic_vector(31 downto 0);
	  output : out std_logic_vector(31 downto 0));
end entity lr;

architecture Dataflow of lr is
begin

	output <=
end architecture Dataflow;